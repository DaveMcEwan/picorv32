// This is free and unencumbered software released into the public domain.
//
// Anyone is free to copy, modify, publish, use, compile, sell, or
// distribute this software, either in source code form or as a compiled
// binary, for any purpose, commercial or non-commercial, and by any
// means.

`timescale 1 ns / 1 ps

`ifndef VERILATOR
module testbench #(
  parameter AXI_TEST = 0,
  parameter VERBOSE = 0
);
  reg clk = 1;
  reg resetn = 0;
  wire trap;

  always #5 clk = ~clk;

  initial begin
    repeat (100) @(posedge clk);
    resetn <= 1;
  end

  integer dumplevel;
  initial begin
    if ($test$plusargs("vcd")) begin
      $dumpfile("testbench.vcd");
      if (!$value$plusargs("dumplevel=%d", dumplevel))
        dumplevel = 0;
      if ($test$plusargs("eva")) begin
        $dumpvars(dumplevel, evmon);
        $dumpoff();
      end
      else
        $dumpvars(dumplevel, testbench);
    end
    repeat (1000000) @(posedge clk);
    $display("TIMEOUT");
    $finish;
  end

  wire trace_valid;
  wire [35:0] trace_data;
  integer trace_file;

  initial begin
    if ($test$plusargs("trace")) begin
      trace_file = $fopen("testbench.trace", "w");
      repeat (10) @(posedge clk);
      while (!trap) begin
        @(posedge clk);
        if (trace_valid)
          $fwrite(trace_file, "%x\n", trace_data);
      end
      $fclose(trace_file);
      $display("Finished writing testbench.trace.");
    end
  end

  picorv32_wrapper #(
    .AXI_TEST (AXI_TEST),
    .VERBOSE  (VERBOSE)
  ) top (
    .clk(clk),
    .resetn(resetn),
    .trap(trap),
    .trace_valid(trace_valid),
    .trace_data(trace_data)
  );

  riscvsys_monitor evmon ( // {{{
    .instr_lui          (top.uut.picorv32_core.instr_lui         ),
    .instr_auipc        (top.uut.picorv32_core.instr_auipc       ),
    .instr_jal          (top.uut.picorv32_core.instr_jal         ),
    .instr_jalr         (top.uut.picorv32_core.instr_jalr        ),
    .instr_beq          (top.uut.picorv32_core.instr_beq         ),
    .instr_bne          (top.uut.picorv32_core.instr_bne         ),
    .instr_blt          (top.uut.picorv32_core.instr_blt         ),
    .instr_bge          (top.uut.picorv32_core.instr_bge         ),
    .instr_bltu         (top.uut.picorv32_core.instr_bltu        ),
    .instr_bgeu         (top.uut.picorv32_core.instr_bgeu        ),
    .instr_lb           (top.uut.picorv32_core.instr_lb          ),
    .instr_lh           (top.uut.picorv32_core.instr_lh          ),
    .instr_lw           (top.uut.picorv32_core.instr_lw          ),
    .instr_lbu          (top.uut.picorv32_core.instr_lbu         ),
    .instr_lhu          (top.uut.picorv32_core.instr_lhu         ),
    .instr_sb           (top.uut.picorv32_core.instr_sb          ),
    .instr_sh           (top.uut.picorv32_core.instr_sh          ),
    .instr_sw           (top.uut.picorv32_core.instr_sw          ),
    .instr_addi         (top.uut.picorv32_core.instr_addi        ),
    .instr_slti         (top.uut.picorv32_core.instr_slti        ),
    .instr_sltiu        (top.uut.picorv32_core.instr_sltiu       ),
    .instr_xori         (top.uut.picorv32_core.instr_xori        ),
    .instr_ori          (top.uut.picorv32_core.instr_ori         ),
    .instr_andi         (top.uut.picorv32_core.instr_andi        ),
    .instr_slli         (top.uut.picorv32_core.instr_slli        ),
    .instr_srli         (top.uut.picorv32_core.instr_srli        ),
    .instr_srai         (top.uut.picorv32_core.instr_srai        ),
    .instr_add          (top.uut.picorv32_core.instr_add         ),
    .instr_sub          (top.uut.picorv32_core.instr_sub         ),
    .instr_sll          (top.uut.picorv32_core.instr_sll         ),
    .instr_slt          (top.uut.picorv32_core.instr_slt         ),
    .instr_sltu         (top.uut.picorv32_core.instr_sltu        ),
    .instr_xor          (top.uut.picorv32_core.instr_xor         ),
    .instr_srl          (top.uut.picorv32_core.instr_srl         ),
    .instr_sra          (top.uut.picorv32_core.instr_sra         ),
    .instr_or           (top.uut.picorv32_core.instr_or          ),
    .instr_and          (top.uut.picorv32_core.instr_and         ),
    .instr_rdcycle      (top.uut.picorv32_core.instr_rdcycle     ),
    .instr_rdcycleh     (top.uut.picorv32_core.instr_rdcycleh    ),
    .instr_rdinstr      (top.uut.picorv32_core.instr_rdinstr     ),
    .instr_rdinstrh     (top.uut.picorv32_core.instr_rdinstrh    ),
    .instr_ecall_ebreak (top.uut.picorv32_core.instr_ecall_ebreak),
    .instr_getq         (top.uut.picorv32_core.instr_getq        ),
    .instr_setq         (top.uut.picorv32_core.instr_setq        ),
    .instr_retirq       (top.uut.picorv32_core.instr_retirq      ),
    .instr_maskirq      (top.uut.picorv32_core.instr_maskirq     ),
    .instr_waitirq      (top.uut.picorv32_core.instr_waitirq     ),
    .instr_timer        (top.uut.picorv32_core.instr_timer       ),
    .instr_trap         (top.uut.picorv32_core.instr_trap        ),
    .dbg_next (top.uut.picorv32_core.dbg_next)
  ); // }}}

endmodule
`endif

module riscvsys_monitor ( // {{{
  input wire instr_lui,
  input wire instr_auipc,
  input wire instr_jal,
  input wire instr_jalr,
  input wire instr_beq,
  input wire instr_bne,
  input wire instr_blt,
  input wire instr_bge,
  input wire instr_bltu,
  input wire instr_bgeu,
  input wire instr_lb,
  input wire instr_lh,
  input wire instr_lw,
  input wire instr_lbu,
  input wire instr_lhu,
  input wire instr_sb,
  input wire instr_sh,
  input wire instr_sw,
  input wire instr_addi,
  input wire instr_slti,
  input wire instr_sltiu,
  input wire instr_xori,
  input wire instr_ori,
  input wire instr_andi,
  input wire instr_slli,
  input wire instr_srli,
  input wire instr_srai,
  input wire instr_add,
  input wire instr_sub,
  input wire instr_sll,
  input wire instr_slt,
  input wire instr_sltu,
  input wire instr_xor,
  input wire instr_srl,
  input wire instr_sra,
  input wire instr_or,
  input wire instr_and,
  input wire instr_rdcycle,
  input wire instr_rdcycleh,
  input wire instr_rdinstr,
  input wire instr_rdinstrh,
  input wire instr_ecall_ebreak,
  input wire instr_getq,
  input wire instr_setq,
  input wire instr_retirq,
  input wire instr_maskirq,
  input wire instr_waitirq,
  input wire instr_timer,
  input wire instr_trap,
  input wire dbg_next
);
  wire next_lui           = dbg_next && instr_lui;
  wire next_auipc         = dbg_next && instr_auipc;
  wire next_jal           = dbg_next && instr_jal;
  wire next_jalr          = dbg_next && instr_jalr;
  wire next_beq           = dbg_next && instr_beq;
  wire next_bne           = dbg_next && instr_bne;
  wire next_blt           = dbg_next && instr_blt;
  wire next_bge           = dbg_next && instr_bge;
  wire next_bltu          = dbg_next && instr_bltu;
  wire next_bgeu          = dbg_next && instr_bgeu;
  wire next_lb            = dbg_next && instr_lb;
  wire next_lh            = dbg_next && instr_lh;
  wire next_lw            = dbg_next && instr_lw;
  wire next_lbu           = dbg_next && instr_lbu;
  wire next_lhu           = dbg_next && instr_lhu;
  wire next_sb            = dbg_next && instr_sb;
  wire next_sh            = dbg_next && instr_sh;
  wire next_sw            = dbg_next && instr_sw;
  wire next_addi          = dbg_next && instr_addi;
  wire next_slti          = dbg_next && instr_slti;
  wire next_sltiu         = dbg_next && instr_sltiu;
  wire next_xori          = dbg_next && instr_xori;
  wire next_ori           = dbg_next && instr_ori;
  wire next_andi          = dbg_next && instr_andi;
  wire next_slli          = dbg_next && instr_slli;
  wire next_srli          = dbg_next && instr_srli;
  wire next_srai          = dbg_next && instr_srai;
  wire next_add           = dbg_next && instr_add;
  wire next_sub           = dbg_next && instr_sub;
  wire next_sll           = dbg_next && instr_sll;
  wire next_slt           = dbg_next && instr_slt;
  wire next_sltu          = dbg_next && instr_sltu;
  wire next_xor           = dbg_next && instr_xor;
  wire next_srl           = dbg_next && instr_srl;
  wire next_sra           = dbg_next && instr_sra;
  wire next_or            = dbg_next && instr_or;
  wire next_and           = dbg_next && instr_and;
  wire next_rdcycle       = dbg_next && instr_rdcycle;
  wire next_rdcycleh      = dbg_next && instr_rdcycleh;
  wire next_rdinstr       = dbg_next && instr_rdinstr;
  wire next_rdinstrh      = dbg_next && instr_rdinstrh;
  wire next_ecall_ebreak  = dbg_next && instr_ecall_ebreak;
  wire next_getq          = dbg_next && instr_getq;
  wire next_setq          = dbg_next && instr_setq;
  wire next_retirq        = dbg_next && instr_retirq;
  wire next_maskirq       = dbg_next && instr_maskirq;
  wire next_waitirq       = dbg_next && instr_waitirq;
  wire next_timer         = dbg_next && instr_timer;
  wire next_trap          = dbg_next && instr_trap;
endmodule // }}}

module picorv32_wrapper #(
  parameter AXI_TEST = 0,
  parameter VERBOSE = 0
) (
  input clk,
  input resetn,
  output trap,
  output trace_valid,
  output [35:0] trace_data
);
  wire tests_passed;
  reg [31:0] irq;

  always @* begin
    irq = 0;
    irq[4] = &uut.picorv32_core.count_cycle[12:0];
    irq[5] = &uut.picorv32_core.count_cycle[15:0];
  end

  wire        mem_axi_awvalid;
  wire        mem_axi_awready;
  wire [31:0] mem_axi_awaddr;
  wire [ 2:0] mem_axi_awprot;

  wire        mem_axi_wvalid;
  wire        mem_axi_wready;
  wire [31:0] mem_axi_wdata;
  wire [ 3:0] mem_axi_wstrb;

  wire        mem_axi_bvalid;
  wire        mem_axi_bready;

  wire        mem_axi_arvalid;
  wire        mem_axi_arready;
  wire [31:0] mem_axi_araddr;
  wire [ 2:0] mem_axi_arprot;

  wire        mem_axi_rvalid;
  wire        mem_axi_rready;
  wire [31:0] mem_axi_rdata;

  axi4_memory #(
    .AXI_TEST (AXI_TEST),
    .VERBOSE  (VERBOSE)
  ) mem (
    .clk             (clk             ),
    .mem_axi_awvalid (mem_axi_awvalid ),
    .mem_axi_awready (mem_axi_awready ),
    .mem_axi_awaddr  (mem_axi_awaddr  ),
    .mem_axi_awprot  (mem_axi_awprot  ),

    .mem_axi_wvalid  (mem_axi_wvalid  ),
    .mem_axi_wready  (mem_axi_wready  ),
    .mem_axi_wdata   (mem_axi_wdata   ),
    .mem_axi_wstrb   (mem_axi_wstrb   ),

    .mem_axi_bvalid  (mem_axi_bvalid  ),
    .mem_axi_bready  (mem_axi_bready  ),

    .mem_axi_arvalid (mem_axi_arvalid ),
    .mem_axi_arready (mem_axi_arready ),
    .mem_axi_araddr  (mem_axi_araddr  ),
    .mem_axi_arprot  (mem_axi_arprot  ),

    .mem_axi_rvalid  (mem_axi_rvalid  ),
    .mem_axi_rready  (mem_axi_rready  ),
    .mem_axi_rdata   (mem_axi_rdata   ),

    .tests_passed    (tests_passed    )
  );

`ifdef RISCV_FORMAL
  wire        rvfi_valid;
  wire [63:0] rvfi_order;
  wire [31:0] rvfi_insn;
  wire        rvfi_trap;
  wire        rvfi_halt;
  wire        rvfi_intr;
  wire [4:0]  rvfi_rs1_addr;
  wire [4:0]  rvfi_rs2_addr;
  wire [31:0] rvfi_rs1_rdata;
  wire [31:0] rvfi_rs2_rdata;
  wire [4:0]  rvfi_rd_addr;
  wire [31:0] rvfi_rd_wdata;
  wire [31:0] rvfi_pc_rdata;
  wire [31:0] rvfi_pc_wdata;
  wire [31:0] rvfi_mem_addr;
  wire [3:0]  rvfi_mem_rmask;
  wire [3:0]  rvfi_mem_wmask;
  wire [31:0] rvfi_mem_rdata;
  wire [31:0] rvfi_mem_wdata;
`endif

  picorv32_axi #(
`ifndef SYNTH_TEST
`ifdef SP_TEST
    .ENABLE_REGS_DUALPORT(0),
`endif
`ifdef COMPRESSED_ISA
    .COMPRESSED_ISA(1),
`endif
    .ENABLE_MUL(1),
    .ENABLE_DIV(1),
    .ENABLE_IRQ(1),
    .ENABLE_TRACE(1)
`endif
  ) uut (
    .clk            (clk            ),
    .resetn         (resetn         ),
    .trap           (trap           ),
    .mem_axi_awvalid(mem_axi_awvalid),
    .mem_axi_awready(mem_axi_awready),
    .mem_axi_awaddr (mem_axi_awaddr ),
    .mem_axi_awprot (mem_axi_awprot ),
    .mem_axi_wvalid (mem_axi_wvalid ),
    .mem_axi_wready (mem_axi_wready ),
    .mem_axi_wdata  (mem_axi_wdata  ),
    .mem_axi_wstrb  (mem_axi_wstrb  ),
    .mem_axi_bvalid (mem_axi_bvalid ),
    .mem_axi_bready (mem_axi_bready ),
    .mem_axi_arvalid(mem_axi_arvalid),
    .mem_axi_arready(mem_axi_arready),
    .mem_axi_araddr (mem_axi_araddr ),
    .mem_axi_arprot (mem_axi_arprot ),
    .mem_axi_rvalid (mem_axi_rvalid ),
    .mem_axi_rready (mem_axi_rready ),
    .mem_axi_rdata  (mem_axi_rdata  ),
    .irq            (irq            ),
`ifdef RISCV_FORMAL
    .rvfi_valid     (rvfi_valid     ),
    .rvfi_order     (rvfi_order     ),
    .rvfi_insn      (rvfi_insn      ),
    .rvfi_trap      (rvfi_trap      ),
    .rvfi_halt      (rvfi_halt      ),
    .rvfi_intr      (rvfi_intr      ),
    .rvfi_rs1_addr  (rvfi_rs1_addr  ),
    .rvfi_rs2_addr  (rvfi_rs2_addr  ),
    .rvfi_rs1_rdata (rvfi_rs1_rdata ),
    .rvfi_rs2_rdata (rvfi_rs2_rdata ),
    .rvfi_rd_addr   (rvfi_rd_addr   ),
    .rvfi_rd_wdata  (rvfi_rd_wdata  ),
    .rvfi_pc_rdata  (rvfi_pc_rdata  ),
    .rvfi_pc_wdata  (rvfi_pc_wdata  ),
    .rvfi_mem_addr  (rvfi_mem_addr  ),
    .rvfi_mem_rmask (rvfi_mem_rmask ),
    .rvfi_mem_wmask (rvfi_mem_wmask ),
    .rvfi_mem_rdata (rvfi_mem_rdata ),
    .rvfi_mem_wdata (rvfi_mem_wdata ),
`endif
    .trace_valid    (trace_valid    ),
    .trace_data     (trace_data     )
  );

`ifdef RISCV_FORMAL
  picorv32_rvfimon rvfi_monitor (
    .clock          (clk           ),
    .reset          (!resetn       ),
    .rvfi_valid     (rvfi_valid    ),
    .rvfi_order     (rvfi_order    ),
    .rvfi_insn      (rvfi_insn     ),
    .rvfi_trap      (rvfi_trap     ),
    .rvfi_halt      (rvfi_halt     ),
    .rvfi_intr      (rvfi_intr     ),
    .rvfi_rs1_addr  (rvfi_rs1_addr ),
    .rvfi_rs2_addr  (rvfi_rs2_addr ),
    .rvfi_rs1_rdata (rvfi_rs1_rdata),
    .rvfi_rs2_rdata (rvfi_rs2_rdata),
    .rvfi_rd_addr   (rvfi_rd_addr  ),
    .rvfi_rd_wdata  (rvfi_rd_wdata ),
    .rvfi_pc_rdata  (rvfi_pc_rdata ),
    .rvfi_pc_wdata  (rvfi_pc_wdata ),
    .rvfi_mem_addr  (rvfi_mem_addr ),
    .rvfi_mem_rmask (rvfi_mem_rmask),
    .rvfi_mem_wmask (rvfi_mem_wmask),
    .rvfi_mem_rdata (rvfi_mem_rdata),
    .rvfi_mem_wdata (rvfi_mem_wdata)
  );
`endif

  reg [1023:0] firmware_file;
  initial begin
    if (!$value$plusargs("firmware=%s", firmware_file))
      firmware_file = "firmware/firmware.hex";
    $readmemh(firmware_file, mem.memory);
  end

  integer cycle_counter;
  always @(posedge clk) begin
    cycle_counter <= resetn ? cycle_counter + 1 : 0;
    if (resetn && trap) begin
`ifndef VERILATOR
      repeat (10) @(posedge clk);
`endif
      $display("TRAP after %1d clock cycles", cycle_counter);
      if (tests_passed) begin
        $display("ALL TESTS PASSED.");
        $finish;
      end else begin
        $display("ERROR!");
        if ($test$plusargs("noerror"))
          $finish;
        $stop;
      end
    end
  end
endmodule

module axi4_memory #(
  parameter AXI_TEST = 0,
  parameter VERBOSE = 0
) (
  input             clk,
  input             mem_axi_awvalid,
  output reg        mem_axi_awready = 0,
  input [31:0]      mem_axi_awaddr,
  input [ 2:0]      mem_axi_awprot,

  input            mem_axi_wvalid,
  output reg       mem_axi_wready = 0,
  input [31:0]     mem_axi_wdata,
  input [ 3:0]     mem_axi_wstrb,

  output reg       mem_axi_bvalid = 0,
  input            mem_axi_bready,

  input            mem_axi_arvalid,
  output reg       mem_axi_arready = 0,
  input [31:0]     mem_axi_araddr,
  input [ 2:0]     mem_axi_arprot,

  output reg        mem_axi_rvalid = 0,
  input             mem_axi_rready,
  output reg [31:0] mem_axi_rdata,

  output reg tests_passed
);
  reg [31:0]   memory [0:64*1024/4-1] /* verilator public */;
  reg verbose;
  initial verbose = $test$plusargs("verbose") || VERBOSE;

  reg axi_test;
  initial axi_test = $test$plusargs("axi_test") || AXI_TEST;

  initial tests_passed = 0;

  reg [63:0] xorshift64_state = 64'd88172645463325252;

  task xorshift64_next;
    begin
      // see page 4 of Marsaglia, George (July 2003). "Xorshift RNGs". Journal of Statistical Software 8 (14).
      xorshift64_state = xorshift64_state ^ (xorshift64_state << 13);
      xorshift64_state = xorshift64_state ^ (xorshift64_state >>  7);
      xorshift64_state = xorshift64_state ^ (xorshift64_state << 17);
    end
  endtask

  reg [2:0] fast_axi_transaction = ~0;
  reg [4:0] async_axi_transaction = ~0;
  reg [4:0] delay_axi_transaction = 0;

  always @(posedge clk) begin
    if (axi_test) begin
        xorshift64_next;
        {fast_axi_transaction, async_axi_transaction, delay_axi_transaction} <= xorshift64_state;
    end
  end

  reg latched_raddr_en = 0;
  reg latched_waddr_en = 0;
  reg latched_wdata_en = 0;

  reg fast_raddr = 0;
  reg fast_waddr = 0;
  reg fast_wdata = 0;

  reg [31:0] latched_raddr;
  reg [31:0] latched_waddr;
  reg [31:0] latched_wdata;
  reg [ 3:0] latched_wstrb;
  reg        latched_rinsn;

  task handle_axi_arvalid; begin
    mem_axi_arready <= 1;
    latched_raddr = mem_axi_araddr;
    latched_rinsn = mem_axi_arprot[2];
    latched_raddr_en = 1;
    fast_raddr <= 1;
  end endtask

  task handle_axi_awvalid; begin
    mem_axi_awready <= 1;
    latched_waddr = mem_axi_awaddr;
    latched_waddr_en = 1;
    fast_waddr <= 1;
  end endtask

  task handle_axi_wvalid; begin
    mem_axi_wready <= 1;
    latched_wdata = mem_axi_wdata;
    latched_wstrb = mem_axi_wstrb;
    latched_wdata_en = 1;
    fast_wdata <= 1;
  end endtask

  task handle_axi_rvalid; begin
    if (verbose)
      $display("RD: ADDR=%08x DATA=%08x%s", latched_raddr, memory[latched_raddr >> 2], latched_rinsn ? " INSN" : "");
    if (latched_raddr < 64*1024) begin
      mem_axi_rdata <= memory[latched_raddr >> 2];
      mem_axi_rvalid <= 1;
      latched_raddr_en = 0;
    end else begin
      $display("OUT-OF-BOUNDS MEMORY READ FROM %08x", latched_raddr);
      $finish;
    end
  end endtask

  task handle_axi_bvalid; begin
    if (verbose)
      $display("WR: ADDR=%08x DATA=%08x STRB=%04b", latched_waddr, latched_wdata, latched_wstrb);
    if (latched_waddr < 64*1024) begin
      if (latched_wstrb[0]) memory[latched_waddr >> 2][ 7: 0] <= latched_wdata[ 7: 0];
      if (latched_wstrb[1]) memory[latched_waddr >> 2][15: 8] <= latched_wdata[15: 8];
      if (latched_wstrb[2]) memory[latched_waddr >> 2][23:16] <= latched_wdata[23:16];
      if (latched_wstrb[3]) memory[latched_waddr >> 2][31:24] <= latched_wdata[31:24];
    end else
    if (latched_waddr == 32'h1000_0000) begin
      if (verbose) begin
        if (32 <= latched_wdata && latched_wdata < 128)
          $display("OUT: '%c'", latched_wdata[7:0]);
        else
          $display("OUT: %3d", latched_wdata);
      end else begin
        $write("%c", latched_wdata[7:0]);
`ifndef VERILATOR
        $fflush();
`endif
      end
    end else
    if (latched_waddr == 32'h2000_0000) begin
      if (latched_wdata == 123456789)
        tests_passed = 1;
      else if (latched_wdata == 32'hcafebabe)
        $dumpon();
    end else begin
      $display("OUT-OF-BOUNDS MEMORY WRITE TO %08x", latched_waddr);
      $finish;
    end
    mem_axi_bvalid <= 1;
    latched_waddr_en = 0;
    latched_wdata_en = 0;
  end endtask

  always @(negedge clk) begin
    if (mem_axi_arvalid && !(latched_raddr_en || fast_raddr) && async_axi_transaction[0]) handle_axi_arvalid;
    if (mem_axi_awvalid && !(latched_waddr_en || fast_waddr) && async_axi_transaction[1]) handle_axi_awvalid;
    if (mem_axi_wvalid  && !(latched_wdata_en || fast_wdata) && async_axi_transaction[2]) handle_axi_wvalid;
    if (!mem_axi_rvalid && latched_raddr_en && async_axi_transaction[3]) handle_axi_rvalid;
    if (!mem_axi_bvalid && latched_waddr_en && latched_wdata_en && async_axi_transaction[4]) handle_axi_bvalid;
  end

  always @(posedge clk) begin
    mem_axi_arready <= 0;
    mem_axi_awready <= 0;
    mem_axi_wready <= 0;

    fast_raddr <= 0;
    fast_waddr <= 0;
    fast_wdata <= 0;

    if (mem_axi_rvalid && mem_axi_rready) begin
      mem_axi_rvalid <= 0;
    end

    if (mem_axi_bvalid && mem_axi_bready) begin
      mem_axi_bvalid <= 0;
    end

    if (mem_axi_arvalid && mem_axi_arready && !fast_raddr) begin
      latched_raddr = mem_axi_araddr;
      latched_rinsn = mem_axi_arprot[2];
      latched_raddr_en = 1;
    end

    if (mem_axi_awvalid && mem_axi_awready && !fast_waddr) begin
      latched_waddr = mem_axi_awaddr;
      latched_waddr_en = 1;
    end

    if (mem_axi_wvalid && mem_axi_wready && !fast_wdata) begin
      latched_wdata = mem_axi_wdata;
      latched_wstrb = mem_axi_wstrb;
      latched_wdata_en = 1;
    end

    if (mem_axi_arvalid && !(latched_raddr_en || fast_raddr) && !delay_axi_transaction[0]) handle_axi_arvalid;
    if (mem_axi_awvalid && !(latched_waddr_en || fast_waddr) && !delay_axi_transaction[1]) handle_axi_awvalid;
    if (mem_axi_wvalid  && !(latched_wdata_en || fast_wdata) && !delay_axi_transaction[2]) handle_axi_wvalid;

    if (!mem_axi_rvalid && latched_raddr_en && !delay_axi_transaction[3]) handle_axi_rvalid;
    if (!mem_axi_bvalid && latched_waddr_en && latched_wdata_en && !delay_axi_transaction[4]) handle_axi_bvalid;
  end
endmodule
